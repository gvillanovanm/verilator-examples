module helloworld_eg1;
    initial begin 
        $display("Hello World"); 
        $finish; 
    end
endmodule
